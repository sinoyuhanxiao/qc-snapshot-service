PG_HOST=10.10.60.212
PG_PORT=5432
PG_DBNAME=mes_prod
PG_USER=postgres
PG_PASSWORD=postgres
MONGO_URI=mongodb://admin:snow123456@10.10.60.212:27017/dev-mes-qc?authSource=admin